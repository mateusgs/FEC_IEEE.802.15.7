library IEEE;
use IEEE.STD_LOGIC_1164.all;

package VLC_PHY_FEC_CONSTANTS is

	type INT_ARRAY is array (integer range <>) of integer;
	constant fec_frame: INT_ARRAY(0 to 1022) := (12, 14, 6, 38, 56, 24, 39, 63, 43, 0, 56, 2, 47, 11, 51, 52, 48, 54, 57, 39, 0, 61, 54, 16, 47, 47, 13, 39, 15, 43, 62, 57, 23, 56, 40, 10, 47, 5, 19, 45, 37, 61, 6, 59, 3, 53, 11, 51, 52, 59, 1, 13, 17, 19, 60, 29, 21, 23, 53, 37, 26, 54, 26, 9, 22, 61, 24, 11, 14, 53, 17, 26, 50, 30, 23, 19, 0, 36, 25, 9, 42, 61, 35, 12, 31, 0, 3, 43, 24, 32, 39, 10, 14, 7, 14, 38, 62, 43, 11, 50, 43, 43, 15, 46, 8, 51, 33, 15, 50, 7, 19, 24, 59, 54, 54, 42, 48, 36, 37, 11, 17, 4, 50, 42, 62, 1, 26, 49, 44, 12, 31, 28, 12, 37, 22, 49, 12, 52, 20, 13, 38, 63, 38, 50, 20, 56, 2, 20, 9, 45, 53, 62, 25, 24, 25, 22, 13, 63, 54, 37, 14, 58, 31, 31, 16, 6, 32, 22, 5, 42, 63, 37, 28, 51, 57, 51, 56, 51, 11, 8, 24, 19, 8, 4, 50, 29, 50, 41, 19, 11, 39, 3, 61, 24, 15, 33, 7, 27, 26, 56, 15, 9, 5, 43, 16, 63, 38, 25, 29, 25, 48, 16, 5, 32, 55, 15, 47, 12, 25, 6, 12, 10, 62, 55, 41, 45, 15, 52, 4, 34, 1, 10, 0, 9, 35, 46, 14, 42, 24, 55, 42, 37, 27, 51, 61, 60, 44, 41, 45, 34, 26, 51, 36, 5, 3, 25, 53, 22, 31, 46, 11, 33, 12, 49, 17, 63, 20, 59, 41, 5, 23, 31, 28, 52, 10, 25, 14, 3, 44, 48, 50, 54, 4, 55, 40, 15, 52, 25, 1, 30, 2, 0, 56, 55, 60, 57, 13, 18, 55, 39, 9, 29, 49, 33, 6, 57, 15, 14, 41, 63, 56, 60, 33, 25, 40, 6, 28, 15, 5, 32, 20, 60, 17, 39, 47, 12, 30, 3, 31, 53, 12, 45, 18, 3, 27, 51, 45, 33, 5, 41, 57, 55, 45, 9, 31, 24, 22, 48, 31, 28, 49, 4, 33, 32, 28, 46, 39, 27, 42, 43, 24, 22, 24, 20, 43, 9, 53, 29, 29, 41, 31, 18, 43, 34, 50, 26, 35, 54, 36, 30, 12, 32, 16, 42, 8, 37, 63, 25, 26, 51, 35, 37, 6, 21, 43, 17, 54, 33, 15, 41, 51, 56, 18, 41, 7, 16, 43, 34, 40, 27, 23, 29, 44, 60, 9, 3, 31, 47, 26, 34, 43, 21, 61, 58, 13, 35, 39, 28, 24, 8, 26, 37, 29, 14, 1, 31, 10, 38, 55, 17, 49, 46, 15, 60, 7, 0, 62, 50, 9, 46, 32, 56, 31, 15, 2, 16, 50, 51, 10, 61, 38, 54, 25, 4, 19, 63, 22, 38, 52, 61, 60, 42, 29, 35, 32, 24, 41, 56, 36, 36, 18, 29, 42, 6, 52, 24, 56, 40, 54, 41, 31, 34, 16, 37, 38, 7, 11, 26, 52, 35, 29, 10, 6, 13, 8, 41, 26, 2, 7, 46, 18, 31, 21, 27, 20, 46, 23, 26, 61, 15, 9, 63, 4, 42, 30, 59, 29, 25, 31, 29, 51, 12, 26, 43, 9, 8, 24, 20, 3, 40, 11, 8, 3, 31, 0, 62, 34, 57, 6, 13, 29, 11, 41, 10, 35, 54, 21, 57, 41, 61, 6, 54, 16, 0, 25, 31, 57, 54, 17, 23, 47, 26, 26, 53, 8, 9, 35, 7, 13, 52, 4, 36, 57, 63, 20, 46, 44, 53, 10, 49, 59, 30, 30, 32, 21, 27, 32, 4, 63, 26, 0, 15, 40, 29, 30, 33, 40, 50, 45, 42, 42, 27, 24, 17, 23, 43, 16, 23, 31, 13, 25, 63, 33, 24, 48, 20, 27, 21, 44, 58, 31, 15, 12, 39, 36, 55, 44, 52, 53, 43, 37, 48, 20, 26, 29, 40, 31, 57, 61, 44, 12, 61, 46, 22, 0, 34, 1, 28, 18, 32, 5, 16, 48, 12, 14, 27, 36, 62, 16, 52, 47, 45, 35, 22, 18, 55, 59, 53, 5, 25, 25, 53, 35, 19, 39, 19, 51, 6, 11, 8, 36, 59, 61, 3, 25, 60, 49, 22, 51, 62, 42, 38, 11, 57, 51, 41, 46, 3, 52, 13, 8, 59, 0, 12, 24, 50, 62, 2, 60, 4, 16, 31, 15, 17, 40, 5, 19, 49, 31, 11, 36, 24, 54, 27, 25, 17, 34, 57, 7, 27, 37, 12, 50, 34, 38, 4, 27, 0, 14, 13, 25, 36, 35, 19, 42, 23, 56, 51, 13, 6, 49, 35, 4, 40, 22, 41, 32, 43, 39, 42, 35, 9, 55, 10, 15, 45, 39, 60, 29, 27, 9, 9, 60, 2, 17, 22, 59, 43, 40, 62, 26, 30, 55, 34, 2, 29, 18, 45, 8, 36, 55, 45, 32, 7, 32, 27, 5, 37, 34, 24, 28, 4, 11, 30, 63, 43, 52, 16, 38, 45, 61, 16, 61, 10, 3, 7, 49, 22, 20, 8, 10, 29, 17, 27, 13, 25, 40, 22, 7, 55, 42, 45, 54, 53, 26, 4, 32, 27, 39, 63, 11, 23, 22, 59, 36, 50, 12, 14, 3, 21, 10, 63, 27, 10, 21, 23, 25, 32, 54, 11, 11, 21, 59, 30, 59, 58, 61, 22, 14, 61, 8, 45, 10, 0, 2, 50, 39, 61, 23, 4, 0, 15, 44, 63, 57, 2, 40, 31, 13, 5, 28, 16, 0, 60, 36, 44, 7, 60, 29, 52, 50, 35, 44, 63, 45, 56, 22, 39, 46, 57, 39, 7, 19, 54, 53, 32, 42, 11, 48, 1, 8, 1, 2, 11, 15, 26, 18, 18, 44, 45, 25, 10, 24, 38, 47, 0, 14, 6, 33, 26, 16, 30, 16, 46, 19, 10, 1, 22, 29, 47, 39, 27, 40, 59, 29, 27, 15, 33, 58, 21, 57, 42, 60, 38, 26, 27, 39, 16, 18, 36, 27, 26, 33, 56, 1, 13, 63, 49, 6, 11, 17, 39, 42, 44, 8, 14, 17, 1, 30, 37, 41, 9, 3, 6, 1, 13, 30, 21, 29, 45, 48, 37, 42, 41, 9, 36, 62, 39, 38, 4, 56, 9, 26);
end package VLC_PHY_FEC_CONSTANTS;

